// ft232h_avalon_sys.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module ft232h_avalon_sys (
		input  wire        clk_clk,                                    //              clk.clk
		input  wire        clk_0_clk,                                  //            clk_0.clk
		output wire        ddr3_pll_sharing_pll_mem_clk,               // ddr3_pll_sharing.pll_mem_clk
		output wire        ddr3_pll_sharing_pll_write_clk,             //                 .pll_write_clk
		output wire        ddr3_pll_sharing_pll_locked,                //                 .pll_locked
		output wire        ddr3_pll_sharing_pll_write_clk_pre_phy_clk, //                 .pll_write_clk_pre_phy_clk
		output wire        ddr3_pll_sharing_pll_addr_cmd_clk,          //                 .pll_addr_cmd_clk
		output wire        ddr3_pll_sharing_pll_avl_clk,               //                 .pll_avl_clk
		output wire        ddr3_pll_sharing_pll_config_clk,            //                 .pll_config_clk
		output wire        ddr3_pll_sharing_pll_mem_phy_clk,           //                 .pll_mem_phy_clk
		output wire        ddr3_pll_sharing_afi_phy_clk,               //                 .afi_phy_clk
		output wire        ddr3_pll_sharing_pll_avl_phy_clk,           //                 .pll_avl_phy_clk
		output wire        ddr3_status_local_init_done,                //      ddr3_status.local_init_done
		output wire        ddr3_status_local_cal_success,              //                 .local_cal_success
		output wire        ddr3_status_local_cal_fail,                 //                 .local_cal_fail
		inout  wire [7:0]  ft232_usb_usb_data,                         //        ft232_usb.usb_data
		output wire        ft232_usb_usb_oe_n,                         //                 .usb_oe_n
		output wire        ft232_usb_usb_rd_n,                         //                 .usb_rd_n
		input  wire        ft232_usb_usb_rxf_n,                        //                 .usb_rxf_n
		output wire        ft232_usb_usb_siwu,                         //                 .usb_siwu
		input  wire        ft232_usb_usb_txe_n,                        //                 .usb_txe_n
		output wire        ft232_usb_usb_wr_n,                         //                 .usb_wr_n
		input  wire        ft232_usb_usb_clock,                        //                 .usb_clock
		output wire [12:0] memory_mem_a,                               //           memory.mem_a
		output wire [2:0]  memory_mem_ba,                              //                 .mem_ba
		output wire [0:0]  memory_mem_ck,                              //                 .mem_ck
		output wire [0:0]  memory_mem_ck_n,                            //                 .mem_ck_n
		output wire [0:0]  memory_mem_cke,                             //                 .mem_cke
		output wire [0:0]  memory_mem_cs_n,                            //                 .mem_cs_n
		output wire [1:0]  memory_mem_dm,                              //                 .mem_dm
		output wire [0:0]  memory_mem_ras_n,                           //                 .mem_ras_n
		output wire [0:0]  memory_mem_cas_n,                           //                 .mem_cas_n
		output wire [0:0]  memory_mem_we_n,                            //                 .mem_we_n
		output wire        memory_mem_reset_n,                         //                 .mem_reset_n
		inout  wire [15:0] memory_mem_dq,                              //                 .mem_dq
		inout  wire [1:0]  memory_mem_dqs,                             //                 .mem_dqs
		inout  wire [1:0]  memory_mem_dqs_n,                           //                 .mem_dqs_n
		output wire [0:0]  memory_mem_odt,                             //                 .mem_odt
		input  wire        oct_rzqin,                                  //              oct.rzqin
		input  wire        reset_reset_n                               //            reset.reset_n
	);

	wire         ddr3_afi_clk_clk;                                          // ddr3:afi_clk -> [ddr3:mp_cmd_clk_0_clk, ddr3:mp_rfifo_clk_0_clk, ddr3:mp_wfifo_clk_0_clk, mm_interconnect_1:ddr3_afi_clk_clk, rst_controller_001:clk]
	wire         pll_outclk0_clk;                                           // pll:outclk_0 -> [cpu:clk, dma:clk, dma_ram:clk, ft232:clk, irq_mapper:clk, jtag_uart:clk, mm_interconnect_0:pll_outclk0_clk, mm_interconnect_1:pll_outclk0_clk, mm_interconnect_2:pll_outclk0_clk, mm_interconnect_3:pll_outclk0_clk, ram:clk, rst_controller:clk, sysid:clock, usb_dma:clk]
	wire         ddr3_afi_reset_reset;                                      // ddr3:afi_reset_n -> [ddr3:mp_cmd_reset_n_0_reset_n, ddr3:mp_rfifo_reset_n_0_reset_n, ddr3:mp_wfifo_reset_n_0_reset_n, rst_controller_001:reset_in0]
	wire         cpu_debug_reset_request_reset;                             // cpu:debug_reset_request -> reset:reset_in1
	wire         reset_reset_out_reset;                                     // reset:reset_out -> [ddr3:global_reset_n, ddr3:soft_reset_n, pll:rst, rst_controller:reset_in0]
	wire  [31:0] cpu_data_master_readdata;                                  // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                               // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                               // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [17:0] cpu_data_master_address;                                   // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                      // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_readdatavalid;                             // mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire         cpu_data_master_write;                                     // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                 // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                           // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [17:0] cpu_instruction_master_address;                            // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                               // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                      // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_0_usb_dma_control_port_slave_chipselect;   // mm_interconnect_0:usb_dma_control_port_slave_chipselect -> usb_dma:dma_ctl_chipselect
	wire  [26:0] mm_interconnect_0_usb_dma_control_port_slave_readdata;     // usb_dma:dma_ctl_readdata -> mm_interconnect_0:usb_dma_control_port_slave_readdata
	wire   [2:0] mm_interconnect_0_usb_dma_control_port_slave_address;      // mm_interconnect_0:usb_dma_control_port_slave_address -> usb_dma:dma_ctl_address
	wire         mm_interconnect_0_usb_dma_control_port_slave_write;        // mm_interconnect_0:usb_dma_control_port_slave_write -> usb_dma:dma_ctl_write_n
	wire  [26:0] mm_interconnect_0_usb_dma_control_port_slave_writedata;    // mm_interconnect_0:usb_dma_control_port_slave_writedata -> usb_dma:dma_ctl_writedata
	wire         mm_interconnect_0_dma_control_port_slave_chipselect;       // mm_interconnect_0:dma_control_port_slave_chipselect -> dma:dma_ctl_chipselect
	wire  [26:0] mm_interconnect_0_dma_control_port_slave_readdata;         // dma:dma_ctl_readdata -> mm_interconnect_0:dma_control_port_slave_readdata
	wire   [2:0] mm_interconnect_0_dma_control_port_slave_address;          // mm_interconnect_0:dma_control_port_slave_address -> dma:dma_ctl_address
	wire         mm_interconnect_0_dma_control_port_slave_write;            // mm_interconnect_0:dma_control_port_slave_write -> dma:dma_ctl_write_n
	wire  [26:0] mm_interconnect_0_dma_control_port_slave_writedata;        // mm_interconnect_0:dma_control_port_slave_writedata -> dma:dma_ctl_writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;            // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;             // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;            // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;         // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;         // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;             // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;          // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;               // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;           // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire         mm_interconnect_0_dma_ram_s1_chipselect;                   // mm_interconnect_0:dma_ram_s1_chipselect -> dma_ram:chipselect
	wire  [31:0] mm_interconnect_0_dma_ram_s1_readdata;                     // dma_ram:readdata -> mm_interconnect_0:dma_ram_s1_readdata
	wire  [10:0] mm_interconnect_0_dma_ram_s1_address;                      // mm_interconnect_0:dma_ram_s1_address -> dma_ram:address
	wire   [3:0] mm_interconnect_0_dma_ram_s1_byteenable;                   // mm_interconnect_0:dma_ram_s1_byteenable -> dma_ram:byteenable
	wire         mm_interconnect_0_dma_ram_s1_write;                        // mm_interconnect_0:dma_ram_s1_write -> dma_ram:write
	wire  [31:0] mm_interconnect_0_dma_ram_s1_writedata;                    // mm_interconnect_0:dma_ram_s1_writedata -> dma_ram:writedata
	wire         mm_interconnect_0_dma_ram_s1_clken;                        // mm_interconnect_0:dma_ram_s1_clken -> dma_ram:clken
	wire         mm_interconnect_0_ram_s1_chipselect;                       // mm_interconnect_0:ram_s1_chipselect -> ram:chipselect
	wire   [7:0] mm_interconnect_0_ram_s1_readdata;                         // ram:readdata -> mm_interconnect_0:ram_s1_readdata
	wire  [15:0] mm_interconnect_0_ram_s1_address;                          // mm_interconnect_0:ram_s1_address -> ram:address
	wire         mm_interconnect_0_ram_s1_write;                            // mm_interconnect_0:ram_s1_write -> ram:write
	wire   [7:0] mm_interconnect_0_ram_s1_writedata;                        // mm_interconnect_0:ram_s1_writedata -> ram:writedata
	wire         mm_interconnect_0_ram_s1_clken;                            // mm_interconnect_0:ram_s1_clken -> ram:clken
	wire         usb_dma_read_master_chipselect;                            // usb_dma:read_chipselect -> mm_interconnect_1:usb_dma_read_master_chipselect
	wire  [31:0] usb_dma_read_master_readdata;                              // mm_interconnect_1:usb_dma_read_master_readdata -> usb_dma:read_readdata
	wire         usb_dma_read_master_waitrequest;                           // mm_interconnect_1:usb_dma_read_master_waitrequest -> usb_dma:read_waitrequest
	wire  [26:0] usb_dma_read_master_address;                               // usb_dma:read_address -> mm_interconnect_1:usb_dma_read_master_address
	wire         usb_dma_read_master_read;                                  // usb_dma:read_read_n -> mm_interconnect_1:usb_dma_read_master_read
	wire         usb_dma_read_master_readdatavalid;                         // mm_interconnect_1:usb_dma_read_master_readdatavalid -> usb_dma:read_readdatavalid
	wire         dma_write_master_chipselect;                               // dma:write_chipselect -> mm_interconnect_1:dma_write_master_chipselect
	wire         dma_write_master_waitrequest;                              // mm_interconnect_1:dma_write_master_waitrequest -> dma:write_waitrequest
	wire  [26:0] dma_write_master_address;                                  // dma:write_address -> mm_interconnect_1:dma_write_master_address
	wire   [3:0] dma_write_master_byteenable;                               // dma:write_byteenable -> mm_interconnect_1:dma_write_master_byteenable
	wire         dma_write_master_write;                                    // dma:write_write_n -> mm_interconnect_1:dma_write_master_write
	wire  [31:0] dma_write_master_writedata;                                // dma:write_writedata -> mm_interconnect_1:dma_write_master_writedata
	wire         mm_interconnect_1_ddr3_avl_0_beginbursttransfer;           // mm_interconnect_1:ddr3_avl_0_beginbursttransfer -> ddr3:avl_burstbegin_0
	wire  [31:0] mm_interconnect_1_ddr3_avl_0_readdata;                     // ddr3:avl_rdata_0 -> mm_interconnect_1:ddr3_avl_0_readdata
	wire         mm_interconnect_1_ddr3_avl_0_waitrequest;                  // ddr3:avl_ready_0 -> mm_interconnect_1:ddr3_avl_0_waitrequest
	wire  [24:0] mm_interconnect_1_ddr3_avl_0_address;                      // mm_interconnect_1:ddr3_avl_0_address -> ddr3:avl_addr_0
	wire         mm_interconnect_1_ddr3_avl_0_read;                         // mm_interconnect_1:ddr3_avl_0_read -> ddr3:avl_read_req_0
	wire   [3:0] mm_interconnect_1_ddr3_avl_0_byteenable;                   // mm_interconnect_1:ddr3_avl_0_byteenable -> ddr3:avl_be_0
	wire         mm_interconnect_1_ddr3_avl_0_readdatavalid;                // ddr3:avl_rdata_valid_0 -> mm_interconnect_1:ddr3_avl_0_readdatavalid
	wire         mm_interconnect_1_ddr3_avl_0_write;                        // mm_interconnect_1:ddr3_avl_0_write -> ddr3:avl_write_req_0
	wire  [31:0] mm_interconnect_1_ddr3_avl_0_writedata;                    // mm_interconnect_1:ddr3_avl_0_writedata -> ddr3:avl_wdata_0
	wire   [2:0] mm_interconnect_1_ddr3_avl_0_burstcount;                   // mm_interconnect_1:ddr3_avl_0_burstcount -> ddr3:avl_size_0
	wire         dma_read_master_chipselect;                                // dma:read_chipselect -> mm_interconnect_2:dma_read_master_chipselect
	wire  [31:0] dma_read_master_readdata;                                  // mm_interconnect_2:dma_read_master_readdata -> dma:read_readdata
	wire         dma_read_master_waitrequest;                               // mm_interconnect_2:dma_read_master_waitrequest -> dma:read_waitrequest
	wire  [17:0] dma_read_master_address;                                   // dma:read_address -> mm_interconnect_2:dma_read_master_address
	wire         dma_read_master_read;                                      // dma:read_read_n -> mm_interconnect_2:dma_read_master_read
	wire         dma_read_master_readdatavalid;                             // mm_interconnect_2:dma_read_master_readdatavalid -> dma:read_readdatavalid
	wire         mm_interconnect_2_dma_ram_s2_chipselect;                   // mm_interconnect_2:dma_ram_s2_chipselect -> dma_ram:chipselect2
	wire  [31:0] mm_interconnect_2_dma_ram_s2_readdata;                     // dma_ram:readdata2 -> mm_interconnect_2:dma_ram_s2_readdata
	wire  [10:0] mm_interconnect_2_dma_ram_s2_address;                      // mm_interconnect_2:dma_ram_s2_address -> dma_ram:address2
	wire   [3:0] mm_interconnect_2_dma_ram_s2_byteenable;                   // mm_interconnect_2:dma_ram_s2_byteenable -> dma_ram:byteenable2
	wire         mm_interconnect_2_dma_ram_s2_write;                        // mm_interconnect_2:dma_ram_s2_write -> dma_ram:write2
	wire  [31:0] mm_interconnect_2_dma_ram_s2_writedata;                    // mm_interconnect_2:dma_ram_s2_writedata -> dma_ram:writedata2
	wire         mm_interconnect_2_dma_ram_s2_clken;                        // mm_interconnect_2:dma_ram_s2_clken -> dma_ram:clken2
	wire         usb_dma_write_master_chipselect;                           // usb_dma:write_chipselect -> mm_interconnect_3:usb_dma_write_master_chipselect
	wire         usb_dma_write_master_waitrequest;                          // mm_interconnect_3:usb_dma_write_master_waitrequest -> usb_dma:write_waitrequest
	wire   [9:0] usb_dma_write_master_address;                              // usb_dma:write_address -> mm_interconnect_3:usb_dma_write_master_address
	wire   [3:0] usb_dma_write_master_byteenable;                           // usb_dma:write_byteenable -> mm_interconnect_3:usb_dma_write_master_byteenable
	wire         usb_dma_write_master_write;                                // usb_dma:write_write_n -> mm_interconnect_3:usb_dma_write_master_write
	wire  [31:0] usb_dma_write_master_writedata;                            // usb_dma:write_writedata -> mm_interconnect_3:usb_dma_write_master_writedata
	wire  [31:0] mm_interconnect_3_ft232_avalon_readdata;                   // ft232:avalon_readdata -> mm_interconnect_3:ft232_avalon_readdata
	wire         mm_interconnect_3_ft232_avalon_waitrequest;                // ft232:avalon_waitrequest -> mm_interconnect_3:ft232_avalon_waitrequest
	wire   [7:0] mm_interconnect_3_ft232_avalon_address;                    // mm_interconnect_3:ft232_avalon_address -> ft232:avalon_address
	wire         mm_interconnect_3_ft232_avalon_read;                       // mm_interconnect_3:ft232_avalon_read -> ft232:avalon_read
	wire         mm_interconnect_3_ft232_avalon_write;                      // mm_interconnect_3:ft232_avalon_write -> ft232:avalon_write
	wire  [31:0] mm_interconnect_3_ft232_avalon_writedata;                  // mm_interconnect_3:ft232_avalon_writedata -> ft232:avalon_writedata
	wire         irq_mapper_receiver0_irq;                                  // usb_dma:dma_ctl_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // dma:dma_ctl_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                  // ft232:rx_almost_full -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                  // ft232:tx_almost_empty -> irq_mapper:receiver4_irq
	wire  [31:0] cpu_irq_irq;                                               // irq_mapper:sender_irq -> cpu:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [cpu:reset_n, dma:system_reset_n, dma_ram:reset, ft232:rst_n, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, mm_interconnect_1:usb_dma_reset_reset_bridge_in_reset_reset, mm_interconnect_2:dma_reset_reset_bridge_in_reset_reset, mm_interconnect_3:usb_dma_reset_reset_bridge_in_reset_reset, ram:reset, rst_translator:in_reset, sysid:reset_n, usb_dma:system_reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [cpu:reset_req, dma_ram:reset_req, ram:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [mm_interconnect_1:ddr3_avl_0_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_1:ddr3_mp_cmd_reset_n_0_reset_bridge_in_reset_reset]

	ft232h_avalon_sys_cpu cpu (
		.clk                                 (pll_outclk0_clk),                                   //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	ft232h_avalon_sys_ddr3 ddr3 (
		.pll_ref_clk                (clk_0_clk),                                       //        pll_ref_clk.clk
		.global_reset_n             (~reset_reset_out_reset),                          //       global_reset.reset_n
		.soft_reset_n               (~reset_reset_out_reset),                          //         soft_reset.reset_n
		.afi_clk                    (ddr3_afi_clk_clk),                                //            afi_clk.clk
		.afi_half_clk               (),                                                //       afi_half_clk.clk
		.afi_reset_n                (ddr3_afi_reset_reset),                            //          afi_reset.reset_n
		.afi_reset_export_n         (),                                                //   afi_reset_export.reset_n
		.mem_a                      (memory_mem_a),                                    //             memory.mem_a
		.mem_ba                     (memory_mem_ba),                                   //                   .mem_ba
		.mem_ck                     (memory_mem_ck),                                   //                   .mem_ck
		.mem_ck_n                   (memory_mem_ck_n),                                 //                   .mem_ck_n
		.mem_cke                    (memory_mem_cke),                                  //                   .mem_cke
		.mem_cs_n                   (memory_mem_cs_n),                                 //                   .mem_cs_n
		.mem_dm                     (memory_mem_dm),                                   //                   .mem_dm
		.mem_ras_n                  (memory_mem_ras_n),                                //                   .mem_ras_n
		.mem_cas_n                  (memory_mem_cas_n),                                //                   .mem_cas_n
		.mem_we_n                   (memory_mem_we_n),                                 //                   .mem_we_n
		.mem_reset_n                (memory_mem_reset_n),                              //                   .mem_reset_n
		.mem_dq                     (memory_mem_dq),                                   //                   .mem_dq
		.mem_dqs                    (memory_mem_dqs),                                  //                   .mem_dqs
		.mem_dqs_n                  (memory_mem_dqs_n),                                //                   .mem_dqs_n
		.mem_odt                    (memory_mem_odt),                                  //                   .mem_odt
		.avl_ready_0                (mm_interconnect_1_ddr3_avl_0_waitrequest),        //              avl_0.waitrequest_n
		.avl_burstbegin_0           (mm_interconnect_1_ddr3_avl_0_beginbursttransfer), //                   .beginbursttransfer
		.avl_addr_0                 (mm_interconnect_1_ddr3_avl_0_address),            //                   .address
		.avl_rdata_valid_0          (mm_interconnect_1_ddr3_avl_0_readdatavalid),      //                   .readdatavalid
		.avl_rdata_0                (mm_interconnect_1_ddr3_avl_0_readdata),           //                   .readdata
		.avl_wdata_0                (mm_interconnect_1_ddr3_avl_0_writedata),          //                   .writedata
		.avl_be_0                   (mm_interconnect_1_ddr3_avl_0_byteenable),         //                   .byteenable
		.avl_read_req_0             (mm_interconnect_1_ddr3_avl_0_read),               //                   .read
		.avl_write_req_0            (mm_interconnect_1_ddr3_avl_0_write),              //                   .write
		.avl_size_0                 (mm_interconnect_1_ddr3_avl_0_burstcount),         //                   .burstcount
		.mp_cmd_clk_0_clk           (ddr3_afi_clk_clk),                                //       mp_cmd_clk_0.clk
		.mp_cmd_reset_n_0_reset_n   (ddr3_afi_reset_reset),                            //   mp_cmd_reset_n_0.reset_n
		.mp_rfifo_clk_0_clk         (ddr3_afi_clk_clk),                                //     mp_rfifo_clk_0.clk
		.mp_rfifo_reset_n_0_reset_n (ddr3_afi_reset_reset),                            // mp_rfifo_reset_n_0.reset_n
		.mp_wfifo_clk_0_clk         (ddr3_afi_clk_clk),                                //     mp_wfifo_clk_0.clk
		.mp_wfifo_reset_n_0_reset_n (ddr3_afi_reset_reset),                            // mp_wfifo_reset_n_0.reset_n
		.local_init_done            (ddr3_status_local_init_done),                     //             status.local_init_done
		.local_cal_success          (ddr3_status_local_cal_success),                   //                   .local_cal_success
		.local_cal_fail             (ddr3_status_local_cal_fail),                      //                   .local_cal_fail
		.oct_rzqin                  (oct_rzqin),                                       //                oct.rzqin
		.pll_mem_clk                (ddr3_pll_sharing_pll_mem_clk),                    //        pll_sharing.pll_mem_clk
		.pll_write_clk              (ddr3_pll_sharing_pll_write_clk),                  //                   .pll_write_clk
		.pll_locked                 (ddr3_pll_sharing_pll_locked),                     //                   .pll_locked
		.pll_write_clk_pre_phy_clk  (ddr3_pll_sharing_pll_write_clk_pre_phy_clk),      //                   .pll_write_clk_pre_phy_clk
		.pll_addr_cmd_clk           (ddr3_pll_sharing_pll_addr_cmd_clk),               //                   .pll_addr_cmd_clk
		.pll_avl_clk                (ddr3_pll_sharing_pll_avl_clk),                    //                   .pll_avl_clk
		.pll_config_clk             (ddr3_pll_sharing_pll_config_clk),                 //                   .pll_config_clk
		.pll_mem_phy_clk            (ddr3_pll_sharing_pll_mem_phy_clk),                //                   .pll_mem_phy_clk
		.afi_phy_clk                (ddr3_pll_sharing_afi_phy_clk),                    //                   .afi_phy_clk
		.pll_avl_phy_clk            (ddr3_pll_sharing_pll_avl_phy_clk)                 //                   .pll_avl_phy_clk
	);

	ft232h_avalon_sys_dma dma (
		.clk                (pll_outclk0_clk),                                     //                clk.clk
		.system_reset_n     (~rst_controller_reset_out_reset),                     //              reset.reset_n
		.dma_ctl_address    (mm_interconnect_0_dma_control_port_slave_address),    // control_port_slave.address
		.dma_ctl_chipselect (mm_interconnect_0_dma_control_port_slave_chipselect), //                   .chipselect
		.dma_ctl_readdata   (mm_interconnect_0_dma_control_port_slave_readdata),   //                   .readdata
		.dma_ctl_write_n    (~mm_interconnect_0_dma_control_port_slave_write),     //                   .write_n
		.dma_ctl_writedata  (mm_interconnect_0_dma_control_port_slave_writedata),  //                   .writedata
		.dma_ctl_irq        (irq_mapper_receiver1_irq),                            //                irq.irq
		.read_address       (dma_read_master_address),                             //        read_master.address
		.read_chipselect    (dma_read_master_chipselect),                          //                   .chipselect
		.read_read_n        (dma_read_master_read),                                //                   .read_n
		.read_readdata      (dma_read_master_readdata),                            //                   .readdata
		.read_readdatavalid (dma_read_master_readdatavalid),                       //                   .readdatavalid
		.read_waitrequest   (dma_read_master_waitrequest),                         //                   .waitrequest
		.write_address      (dma_write_master_address),                            //       write_master.address
		.write_chipselect   (dma_write_master_chipselect),                         //                   .chipselect
		.write_waitrequest  (dma_write_master_waitrequest),                        //                   .waitrequest
		.write_write_n      (dma_write_master_write),                              //                   .write_n
		.write_writedata    (dma_write_master_writedata),                          //                   .writedata
		.write_byteenable   (dma_write_master_byteenable)                          //                   .byteenable
	);

	ft232h_avalon_sys_dma_ram dma_ram (
		.address     (mm_interconnect_0_dma_ram_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_dma_ram_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_dma_ram_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_dma_ram_s1_write),      //       .write
		.readdata    (mm_interconnect_0_dma_ram_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_dma_ram_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_dma_ram_s1_byteenable), //       .byteenable
		.address2    (mm_interconnect_2_dma_ram_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_2_dma_ram_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_2_dma_ram_s2_clken),      //       .clken
		.write2      (mm_interconnect_2_dma_ram_s2_write),      //       .write
		.readdata2   (mm_interconnect_2_dma_ram_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_2_dma_ram_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_2_dma_ram_s2_byteenable), //       .byteenable
		.clk         (pll_outclk0_clk),                         //   clk1.clk
		.reset       (rst_controller_reset_out_reset),          // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req)       //       .reset_req
	);

	ft232h_avalon #(
		.READ_DATA                 (0),
		.WRITE_DATA                (1),
		.RX_FIFO_COUNTER           (2),
		.TX_FIFO_COUNTER           (3),
		.RX_ALMOST_FULL_THRESHOLD  (4),
		.TX_ALMOST_EMPTY_THRESHOLD (5),
		.CLEAR_IRQ                 (6),
		.CONTROL                   (7)
	) ft232 (
		.clk                (pll_outclk0_clk),                            //  clock.clk
		.avalon_address     (mm_interconnect_3_ft232_avalon_address),     // avalon.address
		.avalon_read        (mm_interconnect_3_ft232_avalon_read),        //       .read
		.avalon_readdata    (mm_interconnect_3_ft232_avalon_readdata),    //       .readdata
		.avalon_waitrequest (mm_interconnect_3_ft232_avalon_waitrequest), //       .waitrequest
		.avalon_write       (mm_interconnect_3_ft232_avalon_write),       //       .write
		.avalon_writedata   (mm_interconnect_3_ft232_avalon_writedata),   //       .writedata
		.data               (ft232_usb_usb_data),                         //    usb.usb_data
		.oe_n               (ft232_usb_usb_oe_n),                         //       .usb_oe_n
		.rd_n               (ft232_usb_usb_rd_n),                         //       .usb_rd_n
		.rxf_n              (ft232_usb_usb_rxf_n),                        //       .usb_rxf_n
		.siwu               (ft232_usb_usb_siwu),                         //       .usb_siwu
		.txe_n              (ft232_usb_usb_txe_n),                        //       .usb_txe_n
		.wr_n               (ft232_usb_usb_wr_n),                         //       .usb_wr_n
		.clock              (ft232_usb_usb_clock),                        //       .usb_clock
		.rst_n              (~rst_controller_reset_out_reset),            //  reset.reset_n
		.tx_almost_empty    (irq_mapper_receiver4_irq),                   // tx_irq.irq
		.rx_almost_full     (irq_mapper_receiver3_irq)                    // rx_irq.irq
	);

	ft232h_avalon_sys_jtag_uart jtag_uart (
		.clk            (pll_outclk0_clk),                                           //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver2_irq)                                   //               irq.irq
	);

	ft232h_avalon_sys_pll pll (
		.refclk   (clk_clk),               //  refclk.clk
		.rst      (reset_reset_out_reset), //   reset.reset
		.outclk_0 (pll_outclk0_clk),       // outclk0.clk
		.locked   ()                       // (terminated)
	);

	ft232h_avalon_sys_ram ram (
		.clk        (pll_outclk0_clk),                     //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)   //       .reset_req
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) reset (
		.reset_in0      (~reset_reset_n),                // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                       //       clk.clk
		.reset_out      (reset_reset_out_reset),         // reset_out.reset
		.reset_req      (),                              // (terminated)
		.reset_req_in0  (1'b0),                          // (terminated)
		.reset_req_in1  (1'b0),                          // (terminated)
		.reset_in2      (1'b0),                          // (terminated)
		.reset_req_in2  (1'b0),                          // (terminated)
		.reset_in3      (1'b0),                          // (terminated)
		.reset_req_in3  (1'b0),                          // (terminated)
		.reset_in4      (1'b0),                          // (terminated)
		.reset_req_in4  (1'b0),                          // (terminated)
		.reset_in5      (1'b0),                          // (terminated)
		.reset_req_in5  (1'b0),                          // (terminated)
		.reset_in6      (1'b0),                          // (terminated)
		.reset_req_in6  (1'b0),                          // (terminated)
		.reset_in7      (1'b0),                          // (terminated)
		.reset_req_in7  (1'b0),                          // (terminated)
		.reset_in8      (1'b0),                          // (terminated)
		.reset_req_in8  (1'b0),                          // (terminated)
		.reset_in9      (1'b0),                          // (terminated)
		.reset_req_in9  (1'b0),                          // (terminated)
		.reset_in10     (1'b0),                          // (terminated)
		.reset_req_in10 (1'b0),                          // (terminated)
		.reset_in11     (1'b0),                          // (terminated)
		.reset_req_in11 (1'b0),                          // (terminated)
		.reset_in12     (1'b0),                          // (terminated)
		.reset_req_in12 (1'b0),                          // (terminated)
		.reset_in13     (1'b0),                          // (terminated)
		.reset_req_in13 (1'b0),                          // (terminated)
		.reset_in14     (1'b0),                          // (terminated)
		.reset_req_in14 (1'b0),                          // (terminated)
		.reset_in15     (1'b0),                          // (terminated)
		.reset_req_in15 (1'b0)                           // (terminated)
	);

	ft232h_avalon_sys_sysid sysid (
		.clock    (pll_outclk0_clk),                                //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	ft232h_avalon_sys_usb_dma usb_dma (
		.clk                (pll_outclk0_clk),                                         //                clk.clk
		.system_reset_n     (~rst_controller_reset_out_reset),                         //              reset.reset_n
		.dma_ctl_address    (mm_interconnect_0_usb_dma_control_port_slave_address),    // control_port_slave.address
		.dma_ctl_chipselect (mm_interconnect_0_usb_dma_control_port_slave_chipselect), //                   .chipselect
		.dma_ctl_readdata   (mm_interconnect_0_usb_dma_control_port_slave_readdata),   //                   .readdata
		.dma_ctl_write_n    (~mm_interconnect_0_usb_dma_control_port_slave_write),     //                   .write_n
		.dma_ctl_writedata  (mm_interconnect_0_usb_dma_control_port_slave_writedata),  //                   .writedata
		.dma_ctl_irq        (irq_mapper_receiver0_irq),                                //                irq.irq
		.read_address       (usb_dma_read_master_address),                             //        read_master.address
		.read_chipselect    (usb_dma_read_master_chipselect),                          //                   .chipselect
		.read_read_n        (usb_dma_read_master_read),                                //                   .read_n
		.read_readdata      (usb_dma_read_master_readdata),                            //                   .readdata
		.read_readdatavalid (usb_dma_read_master_readdatavalid),                       //                   .readdatavalid
		.read_waitrequest   (usb_dma_read_master_waitrequest),                         //                   .waitrequest
		.write_address      (usb_dma_write_master_address),                            //       write_master.address
		.write_chipselect   (usb_dma_write_master_chipselect),                         //                   .chipselect
		.write_waitrequest  (usb_dma_write_master_waitrequest),                        //                   .waitrequest
		.write_write_n      (usb_dma_write_master_write),                              //                   .write_n
		.write_writedata    (usb_dma_write_master_writedata),                          //                   .writedata
		.write_byteenable   (usb_dma_write_master_byteenable)                          //                   .byteenable
	);

	ft232h_avalon_sys_mm_interconnect_0 mm_interconnect_0 (
		.pll_outclk0_clk                         (pll_outclk0_clk),                                           //                     pll_outclk0.clk
		.cpu_reset_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                            // cpu_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                 (cpu_data_master_address),                                   //                 cpu_data_master.address
		.cpu_data_master_waitrequest             (cpu_data_master_waitrequest),                               //                                .waitrequest
		.cpu_data_master_byteenable              (cpu_data_master_byteenable),                                //                                .byteenable
		.cpu_data_master_read                    (cpu_data_master_read),                                      //                                .read
		.cpu_data_master_readdata                (cpu_data_master_readdata),                                  //                                .readdata
		.cpu_data_master_readdatavalid           (cpu_data_master_readdatavalid),                             //                                .readdatavalid
		.cpu_data_master_write                   (cpu_data_master_write),                                     //                                .write
		.cpu_data_master_writedata               (cpu_data_master_writedata),                                 //                                .writedata
		.cpu_data_master_debugaccess             (cpu_data_master_debugaccess),                               //                                .debugaccess
		.cpu_instruction_master_address          (cpu_instruction_master_address),                            //          cpu_instruction_master.address
		.cpu_instruction_master_waitrequest      (cpu_instruction_master_waitrequest),                        //                                .waitrequest
		.cpu_instruction_master_read             (cpu_instruction_master_read),                               //                                .read
		.cpu_instruction_master_readdata         (cpu_instruction_master_readdata),                           //                                .readdata
		.cpu_instruction_master_readdatavalid    (cpu_instruction_master_readdatavalid),                      //                                .readdatavalid
		.cpu_debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),             //             cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),               //                                .write
		.cpu_debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),                //                                .read
		.cpu_debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),            //                                .readdata
		.cpu_debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),           //                                .writedata
		.cpu_debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),          //                                .byteenable
		.cpu_debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),         //                                .waitrequest
		.cpu_debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),         //                                .debugaccess
		.dma_control_port_slave_address          (mm_interconnect_0_dma_control_port_slave_address),          //          dma_control_port_slave.address
		.dma_control_port_slave_write            (mm_interconnect_0_dma_control_port_slave_write),            //                                .write
		.dma_control_port_slave_readdata         (mm_interconnect_0_dma_control_port_slave_readdata),         //                                .readdata
		.dma_control_port_slave_writedata        (mm_interconnect_0_dma_control_port_slave_writedata),        //                                .writedata
		.dma_control_port_slave_chipselect       (mm_interconnect_0_dma_control_port_slave_chipselect),       //                                .chipselect
		.dma_ram_s1_address                      (mm_interconnect_0_dma_ram_s1_address),                      //                      dma_ram_s1.address
		.dma_ram_s1_write                        (mm_interconnect_0_dma_ram_s1_write),                        //                                .write
		.dma_ram_s1_readdata                     (mm_interconnect_0_dma_ram_s1_readdata),                     //                                .readdata
		.dma_ram_s1_writedata                    (mm_interconnect_0_dma_ram_s1_writedata),                    //                                .writedata
		.dma_ram_s1_byteenable                   (mm_interconnect_0_dma_ram_s1_byteenable),                   //                                .byteenable
		.dma_ram_s1_chipselect                   (mm_interconnect_0_dma_ram_s1_chipselect),                   //                                .chipselect
		.dma_ram_s1_clken                        (mm_interconnect_0_dma_ram_s1_clken),                        //                                .clken
		.jtag_uart_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //     jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                .write
		.jtag_uart_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                .read
		.jtag_uart_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                .readdata
		.jtag_uart_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                .chipselect
		.ram_s1_address                          (mm_interconnect_0_ram_s1_address),                          //                          ram_s1.address
		.ram_s1_write                            (mm_interconnect_0_ram_s1_write),                            //                                .write
		.ram_s1_readdata                         (mm_interconnect_0_ram_s1_readdata),                         //                                .readdata
		.ram_s1_writedata                        (mm_interconnect_0_ram_s1_writedata),                        //                                .writedata
		.ram_s1_chipselect                       (mm_interconnect_0_ram_s1_chipselect),                       //                                .chipselect
		.ram_s1_clken                            (mm_interconnect_0_ram_s1_clken),                            //                                .clken
		.sysid_control_slave_address             (mm_interconnect_0_sysid_control_slave_address),             //             sysid_control_slave.address
		.sysid_control_slave_readdata            (mm_interconnect_0_sysid_control_slave_readdata),            //                                .readdata
		.usb_dma_control_port_slave_address      (mm_interconnect_0_usb_dma_control_port_slave_address),      //      usb_dma_control_port_slave.address
		.usb_dma_control_port_slave_write        (mm_interconnect_0_usb_dma_control_port_slave_write),        //                                .write
		.usb_dma_control_port_slave_readdata     (mm_interconnect_0_usb_dma_control_port_slave_readdata),     //                                .readdata
		.usb_dma_control_port_slave_writedata    (mm_interconnect_0_usb_dma_control_port_slave_writedata),    //                                .writedata
		.usb_dma_control_port_slave_chipselect   (mm_interconnect_0_usb_dma_control_port_slave_chipselect)    //                                .chipselect
	);

	ft232h_avalon_sys_mm_interconnect_1 mm_interconnect_1 (
		.ddr3_afi_clk_clk                                        (ddr3_afi_clk_clk),                                //                                      ddr3_afi_clk.clk
		.pll_outclk0_clk                                         (pll_outclk0_clk),                                 //                                       pll_outclk0.clk
		.ddr3_avl_0_translator_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),              // ddr3_avl_0_translator_reset_reset_bridge_in_reset.reset
		.ddr3_mp_cmd_reset_n_0_reset_bridge_in_reset_reset       (rst_controller_001_reset_out_reset),              //       ddr3_mp_cmd_reset_n_0_reset_bridge_in_reset.reset
		.usb_dma_reset_reset_bridge_in_reset_reset               (rst_controller_reset_out_reset),                  //               usb_dma_reset_reset_bridge_in_reset.reset
		.dma_write_master_address                                (dma_write_master_address),                        //                                  dma_write_master.address
		.dma_write_master_waitrequest                            (dma_write_master_waitrequest),                    //                                                  .waitrequest
		.dma_write_master_byteenable                             (dma_write_master_byteenable),                     //                                                  .byteenable
		.dma_write_master_chipselect                             (dma_write_master_chipselect),                     //                                                  .chipselect
		.dma_write_master_write                                  (~dma_write_master_write),                         //                                                  .write
		.dma_write_master_writedata                              (dma_write_master_writedata),                      //                                                  .writedata
		.usb_dma_read_master_address                             (usb_dma_read_master_address),                     //                               usb_dma_read_master.address
		.usb_dma_read_master_waitrequest                         (usb_dma_read_master_waitrequest),                 //                                                  .waitrequest
		.usb_dma_read_master_chipselect                          (usb_dma_read_master_chipselect),                  //                                                  .chipselect
		.usb_dma_read_master_read                                (~usb_dma_read_master_read),                       //                                                  .read
		.usb_dma_read_master_readdata                            (usb_dma_read_master_readdata),                    //                                                  .readdata
		.usb_dma_read_master_readdatavalid                       (usb_dma_read_master_readdatavalid),               //                                                  .readdatavalid
		.ddr3_avl_0_address                                      (mm_interconnect_1_ddr3_avl_0_address),            //                                        ddr3_avl_0.address
		.ddr3_avl_0_write                                        (mm_interconnect_1_ddr3_avl_0_write),              //                                                  .write
		.ddr3_avl_0_read                                         (mm_interconnect_1_ddr3_avl_0_read),               //                                                  .read
		.ddr3_avl_0_readdata                                     (mm_interconnect_1_ddr3_avl_0_readdata),           //                                                  .readdata
		.ddr3_avl_0_writedata                                    (mm_interconnect_1_ddr3_avl_0_writedata),          //                                                  .writedata
		.ddr3_avl_0_beginbursttransfer                           (mm_interconnect_1_ddr3_avl_0_beginbursttransfer), //                                                  .beginbursttransfer
		.ddr3_avl_0_burstcount                                   (mm_interconnect_1_ddr3_avl_0_burstcount),         //                                                  .burstcount
		.ddr3_avl_0_byteenable                                   (mm_interconnect_1_ddr3_avl_0_byteenable),         //                                                  .byteenable
		.ddr3_avl_0_readdatavalid                                (mm_interconnect_1_ddr3_avl_0_readdatavalid),      //                                                  .readdatavalid
		.ddr3_avl_0_waitrequest                                  (~mm_interconnect_1_ddr3_avl_0_waitrequest)        //                                                  .waitrequest
	);

	ft232h_avalon_sys_mm_interconnect_2 mm_interconnect_2 (
		.pll_outclk0_clk                       (pll_outclk0_clk),                         //                     pll_outclk0.clk
		.dma_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),          // dma_reset_reset_bridge_in_reset.reset
		.dma_read_master_address               (dma_read_master_address),                 //                 dma_read_master.address
		.dma_read_master_waitrequest           (dma_read_master_waitrequest),             //                                .waitrequest
		.dma_read_master_chipselect            (dma_read_master_chipselect),              //                                .chipselect
		.dma_read_master_read                  (~dma_read_master_read),                   //                                .read
		.dma_read_master_readdata              (dma_read_master_readdata),                //                                .readdata
		.dma_read_master_readdatavalid         (dma_read_master_readdatavalid),           //                                .readdatavalid
		.dma_ram_s2_address                    (mm_interconnect_2_dma_ram_s2_address),    //                      dma_ram_s2.address
		.dma_ram_s2_write                      (mm_interconnect_2_dma_ram_s2_write),      //                                .write
		.dma_ram_s2_readdata                   (mm_interconnect_2_dma_ram_s2_readdata),   //                                .readdata
		.dma_ram_s2_writedata                  (mm_interconnect_2_dma_ram_s2_writedata),  //                                .writedata
		.dma_ram_s2_byteenable                 (mm_interconnect_2_dma_ram_s2_byteenable), //                                .byteenable
		.dma_ram_s2_chipselect                 (mm_interconnect_2_dma_ram_s2_chipselect), //                                .chipselect
		.dma_ram_s2_clken                      (mm_interconnect_2_dma_ram_s2_clken)       //                                .clken
	);

	ft232h_avalon_sys_mm_interconnect_3 mm_interconnect_3 (
		.pll_outclk0_clk                           (pll_outclk0_clk),                            //                         pll_outclk0.clk
		.usb_dma_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),             // usb_dma_reset_reset_bridge_in_reset.reset
		.usb_dma_write_master_address              (usb_dma_write_master_address),               //                usb_dma_write_master.address
		.usb_dma_write_master_waitrequest          (usb_dma_write_master_waitrequest),           //                                    .waitrequest
		.usb_dma_write_master_byteenable           (usb_dma_write_master_byteenable),            //                                    .byteenable
		.usb_dma_write_master_chipselect           (usb_dma_write_master_chipselect),            //                                    .chipselect
		.usb_dma_write_master_write                (~usb_dma_write_master_write),                //                                    .write
		.usb_dma_write_master_writedata            (usb_dma_write_master_writedata),             //                                    .writedata
		.ft232_avalon_address                      (mm_interconnect_3_ft232_avalon_address),     //                        ft232_avalon.address
		.ft232_avalon_write                        (mm_interconnect_3_ft232_avalon_write),       //                                    .write
		.ft232_avalon_read                         (mm_interconnect_3_ft232_avalon_read),        //                                    .read
		.ft232_avalon_readdata                     (mm_interconnect_3_ft232_avalon_readdata),    //                                    .readdata
		.ft232_avalon_writedata                    (mm_interconnect_3_ft232_avalon_writedata),   //                                    .writedata
		.ft232_avalon_waitrequest                  (mm_interconnect_3_ft232_avalon_waitrequest)  //                                    .waitrequest
	);

	ft232h_avalon_sys_irq_mapper irq_mapper (
		.clk           (pll_outclk0_clk),                //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (reset_reset_out_reset),              // reset_in0.reset
		.clk            (pll_outclk0_clk),                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~ddr3_afi_reset_reset),              // reset_in0.reset
		.clk            (ddr3_afi_clk_clk),                   //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
